ARCHITECTURE rtl OF paddle IS

BEGIN

END rtl;