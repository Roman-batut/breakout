ARCHITECTURE rtl OF display IS
BEGIN

   
END rtl;