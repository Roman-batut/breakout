ARCHITECTURE rtl OF brick IS
   
BEGIN

END rtl;