ARCHITECTURE rtl OF game_ctl IS
    
BEGIN

    
END rtl;